`timescale 1ns / 1ps

module and2 (input logic a, b, output logic c);
    assign c = a & b;
endmodule

//I'm making changes to commit to the testing branch!