`timescale 1ns / 1ps

module signExtend (
        input logic [31:0] x,
        input logic [9:0] opcode,
        output logic [63:0] y
);

        always_comb begin

                

        end

endmodule